//Verilog HDL for "lab3", "TxFIFO" "functional"

// Clear is active low - as per doc spec

module TxFIFO (PSEL, PWRITE, PWDATA, CLEAR_B, PCLK, shf_read_ready, TxData, SSPTXINTR, fifo_empty);
parameter	FIFO_Width = 8,
			FIFO_Depth = 4;
	

input PSEL, PWRITE, CLEAR_B, PCLK;
input [7:0] PWDATA;
input shf_read_ready;


output reg [7:0] TxData;
output SSPTXINTR;
output fifo_empty;



// Control Regs
reg [FIFO_Width-1:0] fifo [0:FIFO_Depth-1];
reg [1:0] fifo_write_ptr = 0; // Try using $clog2 or function l8r
reg [1:0] fifo_read_ptr = 0; // Try using $clog2 or function l8r
//

// Data Regs
reg empty, full;
reg [2:0] count;

reg [7:0] data_out;
//

//	Output Assigns
assign SSPTXINTR = (count == FIFO_Depth);		// Fifo full
assign fifo_empty = (count == 0);				// Fifo empty

//


integer i;
always @ (posedge PCLK) begin
	if(!CLEAR_B)begin // Clear all FIFO entries
		for(i = 0; i < FIFO_Depth; i = i + 1)begin
			fifo[i] <= {FIFO_Width{1'b0}};
		end
		// Control Clear
		fifo_read_ptr <= 0;
		fifo_write_ptr <= 0;
		count <= 3'b000;
		// Data Clear
		data_out <= 8'h00;
	end else begin
		if(PSEL && PWRITE)begin // Write a 8-bit entry in FIFO
			if(!SSPTXINTR) begin
				fifo[fifo_write_ptr] <= PWDATA; // Write data to FIFO
				fifo_write_ptr <= fifo_write_ptr + 1;
				count <= count + 1;	
			end 
//		end else if(PSEL && !PWRITE) begin	// Read a 8-bit entry
		end
		if(!fifo_empty && shf_read_ready && PWRITE)begin
			TxData <= fifo[fifo_read_ptr];
			fifo_read_ptr <= fifo_read_ptr + 1;
			count <= count - 1;
		end
		
	end

end

endmodule
